`timescale 1ns / 1ps
module helloworld();
initial begin
$display("Hello ! \nIts start of verilog programming");
end
endmodule
